module ()
endmodule